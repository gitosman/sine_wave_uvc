package wave_uvc_package;

	import uvm_pkg::*;
	`include "uvm_macros.svh"
	
	`include "wave_uvc_packet.sv"
	`include "wave_uvc_seqs.sv"
	`include "wave_uvc_sequencer.sv"
	`include "wave_uvc_driver.sv"
	`include "wave_uvc_agent.sv"
	`include "wave_uvc_env.sv"

endpackage

