interface wave_uvc_interface;

real wave_out;

endinterface
